
module unsaved (
	clk_clk,
	reset_reset_n,
	parallelport2_0_conduit_end_export,
	parallelport2_1_conduit_end_export);	

	input		clk_clk;
	input		reset_reset_n;
	inout	[7:0]	parallelport2_0_conduit_end_export;
	inout	[7:0]	parallelport2_1_conduit_end_export;
endmodule
